module fetch(
    input wire clk,
    input wire [15:0] pc_in,
    input wire [31:0] ram_data,
    input wire ram_busy, ram_cack, ram_data_ready,
    output reg ram_read,
    output reg [31:0] instr_out,
    output reg [15:0] ram_addr,
    output reg ram_addr_ovr,
    output reg pc_hold,
    input wire flag_boot_mode
);

reg [1:0] state;
reg c_acked;
reg [15:0] prev_pc;

initial  state = 2'b0;
initial ram_read = 1'b0;
initial ram_addr_ovr = 1'b0;
initial pc_hold = 1'b0;
initial instr_out = 32'b0;

always @(negedge clk) begin
    if(~flag_boot_mode) begin
        if(pc_in != prev_pc) begin
            pc_hold <= 1'b1;
        end

        case(state)
            2'b0: begin  // IDLE STATE
                if((pc_in != prev_pc || pc_hold)) begin // if pc change fetch new instr
                    ram_read <= 1'b1;
                    ram_addr_ovr <= 1'b1;
                    ram_addr <= pc_in; // fetch instruction pc pointing to
                    instr_out <= 32'b0; // no-op as hold instr
                    state <= 2'b1; // got to next state
                end
            end
            2'b1: begin // RAM READ STATE
                if(~ram_cack && ~c_acked) begin // ram didn't registered command, retry
                    ram_read <= 1'b1;
                    ram_addr_ovr <= 1'b1;
                    ram_read <= 1'b1;
                end else begin
                    ram_read <= 1'b0;
                    c_acked <= 1'b1;
                    if(ram_data_ready) begin // ram read finished
                        ram_addr_ovr <= 1'b0;
                        ram_read <= 1'b0;
                        c_acked <= 1'b0;
                        pc_hold <= 1'b0;
                        instr_out <= ram_data;
                        state <= 2'b0;
                    end else begin // wait for data ready
                        ram_addr_ovr <= 1'b1;
                    end
                end
            end
        endcase
        prev_pc <= pc_in;
    end
end

endmodule